library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  library work;
  use work.Constants.all;
  use work.BDTTypes.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2DnNodes(0 to nTrees - 1) := ((22, 12, 4, 12, 22, 20, 27, -2, -2, -2, -2, -2, -2, -2, -2),
                (27, 13, 9, 11, 18, 15, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 12, 4, 22, 12, 27, 24, -2, -2, -2, -2, -2, -2, -2, -2),
                (27, 5, 15, 5, 0, 9, 22, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 18, 4, 18, 18, 24, 24, -2, -2, -2, -2, -2, -2, -2, -2),
                (26, 18, 11, 18, 16, 4, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (24, 25, 24, 20, 4, 17, 25, -2, -2, -2, -2, -2, -2, -2, -2),
                (13, 11, 27, 23, 17, 12, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (13, 6, 17, 8, 6, 4, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (27, 12, 9, 12, 22, 7, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (24, 25, 24, 27, 24, 17, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 11, 11, 5, 25, 23, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 19, 18, 9, 18, 4, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (13, 11, 12, 23, 11, 14, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (26, 24, 4, 24, 12, 20, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 6, 16, 16, 26, 12, 26, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 0, 17, 4, 20, 4, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (13, 17, 27, 23, 0, 4, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (22, 12, 14, 18, 14, 0, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 18, 14, 20, 18, 18, 24, -2, -2, -2, -2, -2, -2, -2, -2),
                (24, 14, 17, 4, 24, 11, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (24, 18, 27, 19, 12, 20, 24, -2, -2, -2, -2, -2, -2, -2, -2),
                (13, 6, 27, 14, 6, 18, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 19, 21, 17, 17, 24, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (9, 26, 17, 8, 4, 0, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 23, 27, 11, 0, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (10, 21, 22, 19, 20, 26, 25, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 21, 12, 24, 18, 18, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 5, 11, 0, 0, 23, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 0, 23, 5, 14, 0, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 4, 0, 11, 17, 4, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 23, 11, 11, 25, 25, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 11, 0, 22, 23, 24, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 16, 6, 12, 10, 27, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (9, 16, 14, 12, 6, 4, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (26, 18, 18, 18, 12, 12, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 20, 12, 1, 10, 14, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 8, 0, 1, 23, 7, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 13, 23, 23, 23, 0, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 20, 0, 5, 4, 14, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 27, 26, 15, 15, 4, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 11, 22, 23, 23, 10, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 22, 1, 11, 17, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (24, 12, 8, 14, 11, 22, 24, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 1, 10, 2, 2, 12, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 6, 23, 24, 6, 8, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 23, 23, 17, 20, 17, 23, -2, -2, -2, -2, -2, -2, -2, -2),
                (13, 12, 4, 24, 4, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 10, 12, 17, 20, 13, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 0, 17, 17, 11, 0, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 8, 27, 10, 19, 17, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 1, 18, 1, 2, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 5, 6, 17, 0, 24, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 27, 2, 15, 15, 18, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 1, 24, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 12, 14, 14, 20, 12, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 17, 0, 11, 0, 11, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 16, 17, 17, 0, 7, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (22, 4, 16, 16, 20, 17, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 11, 27, 17, 23, 0, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 18, 22, 23, 24, 23, 27, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 1, 17, 1, 12, 23, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 1, 12, 4, 2, 10, 22, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 26, 1, 1, 17, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 10, 0, 23, 17, 17, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 1, 20, 2, 2, 12, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 11, 11, 0, 23, 23, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 0, 11, 11, 19, 27, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 22, 24, 4, 22, 20, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 11, 17, 27, 0, 0, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 12, 10, 24, 18, 9, 24, -2, -2, -2, -2, -2, -2, -2, -2),
                (22, 15, 4, 17, 20, 10, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 0, 11, 22, 25, 27, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 17, 22, 8, 21, 11, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 11, 10, -2, 5, 16, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 27, 17, 11, 11, 13, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 1, 1, 8, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 1, 2, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (13, 0, 22, 0, 17, 16, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 14, 12, 11, 12, 12, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (24, 12, 24, 14, 18, 12, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 18, 20, 24, 17, 26, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 1, 1, 2, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (10, 16, 16, 17, 10, 22, 24, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 23, 12, 27, 23, 10, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (22, 27, 17, 20, 9, 17, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (13, 12, 4, 1, 1, 22, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 1, 12, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 1, 11, 4, 22, 23, 25, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 0, 22, 14, 22, 15, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 1, 1, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 22, 17, 16, 10, 20, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (10, 12, 10, 22, 6, 17, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 20, 12, 12, 6, 20, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 17, 20, 27, 0, 22, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 23, 23, 17, 17, 5, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (27, 24, 11, 18, 17, 17, 17, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 14, 27, 27, 17, 15, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 1, 1, 24, 22, 2, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 2, 1, 24, 8, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2DnNodes(0 to nTrees - 1) := ((3584, 60, -4196, -68, -484, 76, 36, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, 100, 12, 44, -76, 20, 1300, 0, 0, 0, 0, 0, 0, 0, 0),
                (180, -52, -4060, 276, 36, 36, -860, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, 76, 20, -76, 35636, 4, 5132, 0, 0, 0, 0, 0, 0, 0, 0),
                (180, 60, -3636, -68, 84, 532, 844, 0, 0, 0, 0, 0, 0, 0, 0),
                (172, 76, -68, -92, -3748, -4828, 60, 0, 0, 0, 0, 0, 0, 0, 0),
                (-516, 932, 492, 60, -4564, 196, 1188, 0, 0, 0, 0, 0, 0, 0, 0),
                (92, -52, 28, 36, -44, -84, 12, 0, 0, 0, 0, 0, 0, 0, 0),
                (108, -20, -244, 76, 12, -1612, 76, 0, 0, 0, 0, 0, 0, 0, 0),
                (28, 28, 4, -28, 2188, 132, 1940, 0, 0, 0, 0, 0, 0, 0, 0),
                (-532, 304, 1012, 28, -1060, -140, 84, 0, 0, 0, 0, 0, 0, 0, 0),
                (52, 52, 28, 60, 164, -4, -9516, 0, 0, 0, 0, 0, 0, 0, 0),
                (-516, 212, 484, 4, -1068, -5972, 44, 0, 0, 0, 0, 0, 0, 0, 0),
                (84, -44, -36, 28, 28, 84, -12, 0, 0, 0, 0, 0, 0, 0, 0),
                (1188, 508, -3812, -500, 4, 68, 576, 0, 0, 0, 0, 0, 0, 0, 0),
                (52, -60, -3716, -3772, 1188, -84, 148, 0, 0, 0, 0, 0, 0, 0, 0),
                (-100, -13156, -204, -5892, 132, -2004, -60, 0, 0, 0, 0, 0, 0, 0, 0),
                (76, 20, 44, 12, -12428, -4108, 28, 0, 0, 0, 0, 0, 0, 0, 0),
                (8144, 20, 84, 4, 76, 82036, -628, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, -12, 36, 44, 44, 28, 36, 0, 0, 0, 0, 0, 0, 0, 0),
                (-980, 84, 100, -1244, -1588, 36, 44, 0, 0, 0, 0, 0, 0, 0, 0),
                (1164, -492, 36, 92, -28, 84, 1892, 0, 0, 0, 0, 0, 0, 0, 0),
                (156, -20, 28, 36, 12, 76, 12, 0, 0, 0, 0, 0, 0, 0, 0),
                (1084, 68, 28, -36, -356, 1644, 1300, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, 1820, -1108, 36, -6116, -68500, 1292, 0, 0, 0, 0, 0, 0, 0, 0),
                (316, 300, 36, -44, 12988, 116, 40276, 0, 0, 0, 0, 0, 0, 0, 0),
                (-3428, 20, 8144, 108, 148, 1556, 52, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1100, 28, 12, -1580, -1348, 4, 36, 0, 0, 0, 0, 0, 0, 0, 0),
                (77676, 44, 28, -45388, 8140, -12, 156, 0, 0, 0, 0, 0, 0, 0, 0),
                (-60, -6084, -780, -204, 132, -24340, -60, 0, 0, 0, 0, 0, 0, 0, 0),
                (1116, -5828, 69988, 36, -1364, -4552, 1788, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, 468, 12, 20, 1572, 172, -3436, 0, 0, 0, 0, 0, 0, 0, 0),
                (-88668, -28, 86932, 3584, -12, -1228, 4, 0, 0, 0, 0, 0, 0, 0, 0),
                (28, 1004, 68, -68, 2436, 44, -4652, 0, 0, 0, 0, 0, 0, 0, 0),
                (12, -3676, 84, 92, 20, -996, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (116, 52, 1116, -52, 52, 12, 84, 0, 0, 0, 0, 0, 0, 0, 0),
                (-468, 1740, -20, -9008, 20, 52, -12, 0, 0, 0, 0, 0, 0, 0, 0),
                (724, 36, 54268, -12944, 988, 116, 1572, 0, 0, 0, 0, 0, 0, 0, 0),
                (-996, 108, -84, -564, -164, -10332, 14460, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, 116, 5332, -52, -1892, 132, -4, 0, 0, 0, 0, 0, 0, 0, 0),
                (836, 44, 1664, 12, 28, -4052, 1092, 0, 0, 0, 0, 0, 0, 0, 0),
                (-81036, -20, 8872, 1236, -4, -1788, 14664, 0, 0, 0, 0, 0, 0, 0, 0),
                (-4652, -1796, -35664, 300, -228, -36888, 8808, 0, 0, 0, 0, 0, 0, 0, 0),
                (1116, -900, 84, 2012, -36, 4568, 1452, 0, 0, 0, 0, 0, 0, 0, 0),
                (148, 35288, 516, 21680, 36896, -116, -268, 0, 0, 0, 0, 0, 0, 0, 0),
                (1372, -28, 1068, -28, 4, 76, 2124, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1388, -1508, -1164, -1876, 2404, -28, 28, 0, 0, 0, 0, 0, 0, 0, 0),
                (124, 548, -1092, -1148, -4052, -3660, -1308, 0, 0, 0, 0, 0, 0, 0, 0),
                (-6180, -316, -580, -36, 1780, 116, -1036, 0, 0, 0, 0, 0, 0, 0, 0),
                (-68, -5116, -28, -4, -52, 6620, -36, 0, 0, 0, 0, 0, 0, 0, 0),
                (90508, 28, 36, -464, 36, -164, 116, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, 12280, -36, -10224, 5680, -23056, 12, 0, 0, 0, 0, 0, 0, 0, 0),
                (-4604, 132, -84, 220, 7504, -516, 172, 0, 0, 0, 0, 0, 0, 0, 0),
                (51512, 44, 53632, 20, 28, -556, 68920, 0, 0, 0, 0, 0, 0, 0, 0),
                (-42720, -44136, -21992, -52784, 2412, -12192, -21040, 0, 0, 0, 0, 0, 0, 0, 0),
                (4, -12, 36, 36, 68, 12, 124, 0, 0, 0, 0, 0, 0, 0, 0),
                (76, 20, 9644, 12, -4868, 36, -4, 0, 0, 0, 0, 0, 0, 0, 0),
                (-956, -972, -780, 84, -15116, 92, 172, 0, 0, 0, 0, 0, 0, 0, 0),
                (3584, -3972, -1060, 316, 140, -124, 116, 0, 0, 0, 0, 0, 0, 0, 0),
                (1236, -196, 36, -156, -84, -17460, -804, 0, 0, 0, 0, 0, 0, 0, 0),
                (60, 508, 3584, -604, 644, 28, 44, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, 16248, 876, -16640, 188, 820, 1956, 0, 0, 0, 0, 0, 0, 0, 0),
                (-988, -13688, 516, -5428, 29512, -556, 10152, 0, 0, 0, 0, 0, 0, 0, 0),
                (-71632, -79464, 116, -77488, -76336, -76, -20, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1612, -252, -90500, -2060, -2108, 244, -2852, 0, 0, 0, 0, 0, 0, 0, 0),
                (28, 29048, 108, 18000, 27616, 108, -84, 0, 0, 0, 0, 0, 0, 0, 0),
                (72084, -28, 76, 5316, 12, 84, 1944, 0, 0, 0, 0, 0, 0, 0, 0),
                (-44, -4188, 28, -12, 100, 28, 108, 0, 0, 0, 0, 0, 0, 0, 0),
                (1220, 3584, 788, -3988, 5068, 2948, -5436, 0, 0, 0, 0, 0, 0, 0, 0),
                (-276, 60, -20, 36, 52, 4604, -20, 0, 0, 0, 0, 0, 0, 0, 0),
                (-2116, -116, -4060, 252, -52, 4, 1412, 0, 0, 0, 0, 0, 0, 0, 0),
                (8972, 12, -5324, -44, 2308, 2436, -516, 0, 0, 0, 0, 0, 0, 0, 0),
                (-28, -4604, 20, 3584, 108, 28, -20636, 0, 0, 0, 0, 0, 0, 0, 0),
                (92868, 1388, 3584, 36, 28, 76, -3588, 0, 0, 0, 0, 0, 0, 0, 0),
                (-4684, -464, -5172, 0, 100, -3556, -2852, 0, 0, 0, 0, 0, 0, -16, -16),
                (-1324, 36, -860, 108, -68, 84, -732, 0, 0, 0, 0, 0, 0, 0, 0),
                (43992, 24096, 45632, 22568, 13736, 132, 56328, 0, 0, 0, 0, 0, 0, 0, 0),
                (-29600, -29704, -43208, -41008, -23496, -26496, -19384, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, 8636, 3584, -8180, 700, 1172, -68, 0, 0, 0, 0, 0, 0, 0, 0),
                (-6236, 148, 44, -44, 556, -44, -6048, 0, 0, 0, 0, 0, 0, 0, 0),
                (-36, -28, 20, 60, 924, -84, 12, 0, 0, 0, 0, 0, 0, 0, 0),
                (-324, -1268, 2284, -956, 12, 2060, 1348, 0, 0, 0, 0, 0, 0, 0, 0),
                (37016, 20816, 38880, 20088, 10280, 33680, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (-3804, -2972, -436, -220, -4332, 3200, -1404, 0, 0, 0, 0, 0, 0, 0, 0),
                (-86404, -100, 1028, 28, -20, -500, 13688, 0, 0, 0, 0, 0, 0, 0, 0),
                (10964, 36, 228, 2380, 4, -116, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (236, 500, -3884, 11112, 12120, 8012, -1244, 0, 0, 0, 0, 0, 0, 0, 0),
                (-8560, -3208, -12888, -25008, -220, -1904, 8328, 0, 0, 0, 0, 0, 0, 0, 0),
                (-796, -6912, 204, -3956, 10152, -1588, 796, 0, 0, 0, 0, 0, 0, 0, 0),
                (-308, -13472, 8144, 68, 3092, 12, 508, 0, 0, 0, 0, 0, 0, 0, 0),
                (72168, 18032, 78208, 18248, 6664, 75088, 76960, 0, 0, 0, 0, 0, 0, 0, 0),
                (-73968, -1772, -1972, -3356, -1788, 2340, -708, 0, 0, 0, 0, 0, 0, 0, 0),
                (-5644, -68, -5340, -1204, 124, 276, -6068, 0, 0, 0, 0, 0, 0, 0, 0),
                (-12, 60, -20, 60, -84, 44, 92, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, 12, 52, 28, -4604, 4484, 5460, 0, 0, 0, 0, 0, 0, 0, 0),
                (72100, -548, 76, -12, -20, 4, 52, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, -1164, -60, -516, -52, 84, -44, 0, 0, 0, 0, 0, 0, 0, 0),
                (-91988, 100, 44, 36, 116, 20, -3020, 0, 0, 0, 0, 0, 0, 0, 0),
                (-828, -10880, -11584, 540, 10152, -5832, -17000, 0, 0, 0, 0, 0, 0, 0, 0),
                (30760, 42352, 31440, 16240, 27032, -2420, 60, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2DnNodes(0 to nTrees - 1) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 13, 7, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2DnNodes(0 to nTrees - 1) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 14, 8, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2DnNodes(0 to nTrees - 1) := ((0, 0, 0, 0, 0, 0, 0, -4, 4, -1, -5, 0, -4, 2, -1),
                (0, 0, 0, 0, 0, 0, 0, 1, -3, -1, 3, -3, -1, 3, 1),
                (0, 0, 0, 0, 0, 0, 0, 1, -4, 2, -2, -2, -3, -3, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 2, -3, 0, -3, -1, 2, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 1, -2, -4, -2, -3, 1, -3),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, -1, -4, -3, 0, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, -4, -3, -2, 0, 1, -1, -3, -1),
                (0, 0, 0, 0, 0, 0, 0, -3, -1, -2, 0, -3, 2, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, -3, -1, 0, -3, -2, 3, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, -1, 2, 1, -3, -2, 0, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, -3, -2, -2, 0, -1, 1, -3, -1),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, -2, 0, -2, 0, 2, -3),
                (0, 0, 0, 0, 0, 0, 0, -2, -3, -2, 0, 0, 1, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -2, -3, 0, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, -2, -4, 1, -1, 2, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, -2, 0, 0, -3, 0, -3, -2),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -3, -2, -1, 1, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, 1, -2, 3),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, -3, 0, -1, 1, -3, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 0, 1, 0, -4, -2, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, 3, -1, 0, 0, -1, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, -2, -1, -1, 0, -4, -2, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, -2, -1, 0, -1, 2, -2, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, -3, 6, -1, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -3, 1, -3),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 0, -3, -1, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, -2, -1, 1, 0, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 8, -3, -2, -1, 0, 0, -3, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, 0, -2, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -3, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, 2, 1, -1, 0, 1, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, -5, -3, -1, 0, -1, 5, -2),
                (0, 0, 0, 0, 0, 0, 0, 1, -2, 0, -1, -1, 3, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, -3, 1, -3, -1, 0, 0, -2, -1),
                (0, 0, 0, 0, 0, 0, 0, -3, -1, -1, 1, -2, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -2, -1, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, -1, -2, 1, -1, 0, -1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -2, 0, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 2, -1, -5, 3, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, -3, 1, 0, 0, 0, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, 1, -21, 9, 3, 0, -3, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 1, 0, 0, -3, -1, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, -2, 0, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, -2, -1, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, -1, 2, -2, -1, 1, -1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -1, -4, 1, 0, -3, 2),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 8, -2, 1, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -1, 0, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, -3, -1, -1, 0, -1, 1, 2, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -3, -1, -1, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, 3, 7, -1, 3, -1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -3, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -3, 4, 1, -2, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, 1, 0, -1, -2, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 0, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 3, 0, -2, -2, 0, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, -3, 1, -3, 5, 2, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, -3, -1, 1, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, -3, -1, 0, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, -2, 0, 0, 0, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 5, -1, -3, 3, 0, 0, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, -4, 0, -4, -3, -1, 1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 3, -1, -3, -2, 1, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, -1, 1, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, 0, -1, 3),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -1, 0, 1, 0, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -2, 0, 2, -1),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -2, -1, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 6, 0, 0, -2, -3, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 1, -2, 2, 1),
                (0, 0, 0, -29, 0, 0, 0, 1, 3, 0, -2, 0, 0, -29, -29),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, 2, 0, -2, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 1, -3, -1, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -3, -1, -3, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, -2, 3, -3, 0, -2, 1, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, 1, -1, 0, 0, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -1, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, 0, 0, 1, -2, 2, -3),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 0, -3, -1, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 1, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, 0, 0, -3, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 1, -1, 7, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 1, 1, 7, -3, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -2, -1, -3, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, 0, -3, 0, 0, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 4, 0, -4, -1, 0, 0, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -4, -2, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, -3, 4, -2, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 5, -1, 1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, -2, 0, -1, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, 0, -1, -2, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 0, 1, -5, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, -2, 0, 0, 0, 1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, 0, 0, 1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 5, 0, -2, 0, -2, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, 6, -2, -1, 0)
                );
    constant parent : intArray2DnNodes(0 to nTrees - 1) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 4, 4, 5, 5, 6, 6, 3, 3),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2DnNodes(0 to nTrees - 1) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2DnLeaves(0 to nTrees - 1) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2DnNodes(0 to nTrees - 1) := to_tyArray2D(value_int);
      constant threshold : txArray2DnNodes(0 to nTrees - 1) := to_txArray2D(threshold_int);
end Arrays0;