library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_misc.all;
  use ieee.numeric_std.all;

  use work.Constants.all;
  use work.BDTTypes.all;
  package Arrays0 is

    constant initPredict : ty := to_ty(0);
    constant feature : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((19, 11, 4, 11, 19, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 11, 4, 11, 19, 19, 21, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 16, 4, 16, 19, 19, 21, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 10, 22, 10, 20, 19, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (21, 22, 21, 4, 4, 15, 22, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 15, 9, 10, 10, 12, 12, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 16, 10, 14, 16, 15, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 6, 17, 6, 23, 11, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (21, 21, 4, 22, 10, 7, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 5, 0, 0, 23, 0, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 23, 16, 16, 19, 16, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 11, 4, 19, 11, 7, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 6, 16, 6, 13, 9, 16, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 10, 10, 0, 9, 4, 21, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 15, 6, 15, 9, 6, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 9, 16, 17, 16, 16, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (21, 4, 4, 23, 19, 13, 23, -2, -2, -2, -2, -2, -2, -2, -2),
                (23, 15, 19, 15, 10, 16, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (18, 17, 4, 10, 6, 9, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 15, 20, 10, 10, 14, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 0, 19, 4, 13, 5, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 6, 11, 8, 16, 19, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (21, 13, 21, 19, 21, 15, 22, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 10, 10, 0, 20, 20, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 0, 15, 4, 10, 20, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 16, 19, 18, 16, 4, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 16, 9, 11, 16, 14, 6, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 18, 16, 16, 16, 9, 23, -2, -2, -2, -2, -2, -2, -2, -2),
                (7, 23, 11, 16, 6, 9, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 1, 18, 2, 1, 11, 23, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 10, 20, 9, 20, 0, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 10, 10, 0, 20, 18, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 4, 17, 19, 19, 20, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 18, 15, 19, 0, 7, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 9, 1, 23, 18, 1, 2, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 14, 0, 15, 15, 5, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 15, 15, 8, 17, 15, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (21, 21, 23, 8, 6, 19, 21, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 13, 16, 16, 17, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 20, 8, 4, 9, 9, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 0, 15, 15, 22, 0, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 16, 17, 15, 18, 4, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 20, 15, 0, 10, 14, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (4, 14, 12, 10, 9, 15, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 11, 9, 11, 16, 14, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 21, 6, 1, 18, 11, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 1, 9, 2, 6, 14, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 15, 19, 4, 13, 0, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 16, 21, 18, 11, 23, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 19, 15, 9, 16, 18, 5, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 4, 8, 23, 8, 21, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 8, 1, 11, 20, 18, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 4, 17, 20, 14, 20, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 21, 9, 21, 11, 14, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 19, 5, 15, 20, 0, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 13, 16, 16, 4, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 1, 1, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 15, 15, 0, 15, 17, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 12, 15, 4, 11, 20, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 20, 0, 18, 15, 13, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (12, 0, 9, 0, 20, 18, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 9, 1, 14, 1, 2, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 14, 17, 10, 9, 1, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 4, 20, 14, 19, 4, 15, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 12, 11, 1, 4, 1, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 1, 19, 2, 2, 15, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 1, 2, 1, 21, -2, -2, -2, -2, -2, -2, -2, -2),
                (21, 14, 9, 15, 23, 14, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 13, 1, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (9, 14, 4, 11, 4, 18, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 1, 11, 2, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 2, 11, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 10, 1, 14, 22, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 15, 15, 0, 12, 20, 22, -2, -2, -2, -2, -2, -2, -2, -2),
                (14, 19, 9, 15, -2, 19, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 10, 0, 20, 15, 20, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 1, 15, 21, 12, 13, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (14, 4, 9, 19, 19, 19, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 21, 21, 4, 8, 14, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (5, 15, 10, 10, 0, 0, 14, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 0, 15, 10, 10, 0, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (8, 21, 14, 11, 21, 16, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (19, 9, 15, 20, 1, 15, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 16, 21, 1, 11, -2, -2, -2, -2, -2, -2, -2, -2),
                (15, 18, 20, 12, 5, 15, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 13, 21, 1, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 0, 20, 10, 20, 10, 19, -2, -2, -2, -2, -2, -2, -2, -2),
                (6, 18, 8, 14, 4, 21, 18, -2, -2, -2, -2, -2, -2, -2, -2),
                (2, 1, 1, 21, 2, 7, 4, -2, -2, -2, -2, -2, -2, -2, -2),
                (16, 1, 4, 2, 2, 21, 21, -2, -2, -2, -2, -2, -2, -2, -2),
                (3, 3, 0, 0, 8, 20, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 14, 20, 0, 15, 0, 10, -2, -2, -2, -2, -2, -2, -2, -2),
                (9, 14, 8, 15, 15, 19, 9, -2, -2, -2, -2, -2, -2, -2, -2),
                (9, 14, 19, 22, 18, 1, 8, -2, -2, -2, -2, -2, -2, -2, -2),
                (1, 2, 2, 4, 16, 16, 1, -2, -2, -2, -2, -2, -2, -2, -2),
                (0, 13, 4, 5, 20, 11, 13, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 8, 1, 21, 9, 23, 21, -2, -2, -2, -2, -2, -2, -2, -2),
                (11, 1, 15, 21, 23, 4, 0, -2, -2, -2, -2, -2, -2, -2, -2),
                (17, 0, 1, 5, 0, 2, 20, -2, -2, -2, -2, -2, -2, -2, -2),
                (20, 15, 15, 9, 0, 0, 15, -2, -2, -2, -2, -2, -2, -2, -2)
                );
    constant threshold_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((3584, 60, -4196, -68, -428, 76, 1300, 0, 0, 0, 0, 0, 0, 0, 0),
                (180, 44, -4060, -52, 172, 7056, -860, 0, 0, 0, 0, 0, 0, 0, 0),
                (3316, 60, -3684, -68, -2004, 7056, 892, 0, 0, 0, 0, 0, 0, 0, 0),
                (100, 44, 924, -52, -52, 10152, -3884, 0, 0, 0, 0, 0, 0, 0, 0),
                (-516, 1444, 500, -3068, -4268, 196, 1444, 0, 0, 0, 0, 0, 0, 0, 0),
                (7056, -188, 1612, -76, -68, 100, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (172, -84, 60, -3668, 76, 52, -4108, 0, 0, 0, 0, 0, 0, 0, 0),
                (92, 12, 800, -12, 172, 28, -1916, 0, 0, 0, 0, 0, 0, 0, 0),
                (1028, -500, -3428, 412, 68, 172, 572, 0, 0, 0, 0, 0, 0, 0, 0),
                (76, -76, 31756, -20388, 1240, 8740, -5748, 0, 0, 0, 0, 0, 0, 0, 0),
                (-5964, 2596, 484, 44, 3316, -508, 44, 0, 0, 0, 0, 0, 0, 0, 0),
                (8144, -36, -1524, -404, 20, 124, -996, 0, 0, 0, 0, 0, 0, 0, 0),
                (108, 4, -76, -20, 36, -1036, 44, 0, 0, 0, 0, 0, 0, 0, 0),
                (-60, -36, -60, 10052, -2596, -3916, -1060, 0, 0, 0, 0, 0, 0, 0, 0),
                (84, 28, 52, -28, -2284, -76, -4572, 0, 0, 0, 0, 0, 0, 0, 0),
                (-476, -636, 12, 2220, -1076, -12, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (1180, -5220, -3092, 2356, 7056, 84, 3572, 0, 0, 0, 0, 0, 0, 0, 0),
                (116, 164, -2148, -188, 60, 92, -2460, 0, 0, 0, 0, 0, 0, 0, 0),
                (2300, 68, -1916, 28, 12, -4, -1124, 0, 0, 0, 0, 0, 0, 0, 0),
                (284, -44, -84, 4, -44, -3916, 25012, 0, 0, 0, 0, 0, 0, 0, 0),
                (-60, -6884, 6164, -5828, 140, 60, -860, 0, 0, 0, 0, 0, 0, 0, 0),
                (140, -20, 76, 68, 980, -1292, -164, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1236, 84, 468, 3584, -1876, -116, 308, 0, 0, 0, 0, 0, 0, 0, 0),
                (72084, -36, 36, 14972, 28, -28, -20, 0, 0, 0, 0, 0, 0, 0, 0),
                (-52, -12156, 36, -5596, -68, 260, 4, 0, 0, 0, 0, 0, 0, 0, 0),
                (-6068, -12, 8144, 52, 4, -3580, -580, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1180, -100, -4076, -52, 84, -3644, 4, 0, 0, 0, 0, 0, 0, 0, 0),
                (-468, 1740, 1124, -516, -1204, -3428, 2420, 0, 0, 0, 0, 0, 0, 0, 0),
                (148, 124, -92, 52, -12, -800, 92, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, -12224, 92, -5320, 11000, -28, 1924, 0, 0, 0, 0, 0, 0, 0, 0),
                (-80420, -76, -28, -92, 1220, -5116, 28, 0, 0, 0, 0, 0, 0, 0, 0),
                (54548, -28, 20, 8500, 12, 1972, -20, 0, 0, 0, 0, 0, 0, 0, 0),
                (1116, -3412, 2220, -2276, 5068, 1012, 1764, 0, 0, 0, 0, 0, 0, 0, 0),
                (-116, 60, -1124, 5260, -12884, 116, -948, 0, 0, 0, 0, 0, 0, 0, 0),
                (8872, -2476, 15560, 3076, 140, -15312, 9376, 0, 0, 0, 0, 0, 0, 0, 0),
                (-60, -4580, -86612, -324, 172, 44, 80820, 0, 0, 0, 0, 0, 0, 0, 0),
                (76, 852, 300, 36, 1964, -292, -2944, 0, 0, 0, 0, 0, 0, 0, 0),
                (1324, -1148, 2876, 84, -20, 3584, 1620, 0, 0, 0, 0, 0, 0, 0, 0),
                (-20, 44, -12, 28, 148, 44, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1372, -708, 28, -3892, 1280, -464, -2892, 0, 0, 0, 0, 0, 0, 0, 0),
                (-276, -15708, -36, -12, 1828, 12524, -28, 0, 0, 0, 0, 0, 0, 0, 0),
                (604, 452, 100, 724, 1756, -3964, 1116, 0, 0, 0, 0, 0, 0, 0, 0),
                (972, -52, 20, -5868, 36, -940, 9844, 0, 0, 0, 0, 0, 0, 0, 0),
                (-6212, -4652, 76, 412, 72, -652, -3756, 0, 0, 0, 0, 0, 0, 0, 0),
                (-436, 84, -4060, -108, 12, -2844, 5276, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1276, -564, 12, 10184, 2948, -868, 84, 0, 0, 0, 0, 0, 0, 0, 0),
                (164, -35616, -2404, -36328, 20, -1076, 124, 0, 0, 0, 0, 0, 0, 0, 0),
                (172, 1372, 3200, -2892, 116, -10788, 4, 0, 0, 0, 0, 0, 0, 0, 0),
                (1196, -20, 796, 76, -12, 2748, -12624, 0, 0, 0, 0, 0, 0, 0, 0),
                (89244, 8980, -260, -548, 508, 2140, 12, 0, 0, 0, 0, 0, 0, 0, 0),
                (5332, -4044, 68, 2380, 68, -724, -1364, 0, 0, 0, 0, 0, 0, 0, 0),
                (748, 28, 12976, -844, 76, 2012, -4004, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1668, -3964, 60, -1772, 3860, -740, -3868, 0, 0, 0, 0, 0, 0, 0, 0),
                (-2060, 68, -4812, -68, -68, -3644, -436, 0, 0, 0, 0, 0, 0, 0, 0),
                (-89732, 3316, -44, 140, -12, -4596, 284, 0, 0, 0, 0, 0, 0, 0, 0),
                (-12, 36, 4, -36, -4260, 68, 36, 0, 0, 0, 0, 0, 0, 0, 0),
                (35256, 20720, 36848, 20424, 10280, 30784, 50360, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1252, -60, -812, 1268, 68, 1700, -2300, 0, 0, 0, 0, 0, 0, 0, 0),
                (-716, 108, 20, -5428, -1284, 484, -69988, 0, 0, 0, 0, 0, 0, 0, 0),
                (52, -44, 6244, 52, -36, 132, -5604, 0, 0, 0, 0, 0, 0, 0, 0),
                (44, 5332, 44, -3556, -12, 2404, -5332, 0, 0, 0, 0, 0, 0, 0, 0),
                (9476, -3516, -8880, -2132, -28048, -2216, 8520, 0, 0, 0, 0, 0, 0, 0, 0),
                (500, -4652, 100, -252, -5172, 6216, 1140, 0, 0, 0, 0, 0, 0, 0, 0),
                (1500, -380, 1204, -268, 7780, -5524, 2124, 0, 0, 0, 0, 0, 0, 0, 0),
                (-580, 544, 12, -6784, -3960, 27800, 60, 0, 0, 0, 0, 0, 0, 0, 0),
                (90668, -70240, 3584, -77016, -19224, -124, -52, 0, 0, 0, 0, 0, 0, 0, 0),
                (-20352, -17960, -33704, -37168, -13960, -12784, 676, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1644, -3500, -3812, 156, 3908, -2724, 5332, 0, 0, 0, 0, 0, 0, 0, 0),
                (-25728, -26152, -40616, 60, -30208, -28, 8776, 0, 0, 0, 0, 0, 0, 0, 0),
                (44, 3316, -5364, -28, -3932, 1804, 1740, 0, 0, 0, 0, 0, 0, 0, 0),
                (17952, 18248, 6520, 12, 11904, 3464, 36744, 0, 0, 0, 0, 0, 0, 0, 0),
                (-8912, -3272, -12888, -10376, -92, -3520, 8776, 0, 0, 0, 0, 0, 0, 0, 0),
                (-60032, -70600, -196, -75904, -3136, 796, -724, 0, 0, 0, 0, 0, 0, 0, 0),
                (-180, 84, 100, 8028, 124, 60, 540, 0, 0, 0, 0, 0, 0, 0, 0),
                (-4564, 348, -5292, 220, 0, -2764, -6180, 0, 0, 0, 0, 0, 0, -16, -16),
                (-70252, -4, 39548, 1364, 4, 580, -4, 0, 0, 0, 0, 0, 0, 0, 0),
                (-996, -13808, 1756, 540, 544, 156, -1476, 0, 0, 0, 0, 0, 0, 0, 0),
                (-260, -4460, -1868, 3316, 2312, 3584, 2200, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1060, -548, -1852, -3924, 76, -1492, 564, 0, 0, 0, 0, 0, 0, 0, 0),
                (52, 20, 92, 20, -4740, 5212, -4172, 0, 0, 0, 0, 0, 0, 0, 0),
                (-68, -9356, -20, -4, -52, 8156, 100, 0, 0, 0, 0, 0, 0, 0, 0),
                (36, -508, 284, 188, 508, -44, 3584, 0, 0, 0, 0, 0, 0, 0, 0),
                (10964, -556, 180, -60, 36936, -148, -9516, 0, 0, 0, 0, 0, 0, 0, 0),
                (-23056, -20872, -35272, -52, 2436, -18832, -12, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1876, 2308, 28, 108, -36, 12, 52, 0, 0, 0, 0, 0, 0, 0, 0),
                (-34608, -32664, -19400, 84, 1180, -7216, -16960, 0, 0, 0, 0, 0, 0, 0, 0),
                (86700, -56044, 100, -12, -748, -100, 3316, 0, 0, 0, 0, 0, 0, 0, 0),
                (-28, 1448, 36, -3756, -3328, -548, 92, 0, 0, 0, 0, 0, 0, 0, 0),
                (48896, 43992, 31816, 1548, 45584, 172, -4004, 0, 0, 0, 0, 0, 0, 0, 0),
                (1380, 73480, -3892, 17952, 78272, 796, 804, 0, 0, 0, 0, 0, 0, 0, 0),
                (-2864, -4480, 29508, -13484, 84, 476, 12, 0, 0, 0, 0, 0, 0, 0, 0),
                (-1380, -972, 76, 11120, -36, 73060, 76, 0, 0, 0, 0, 0, 0, 0, 0),
                (-5068, -3884, 148, 236, 340, -1700, -4364, 0, 0, 0, 0, 0, 0, 0, 0),
                (-708, 332, 6164, 116, 76, 23832, 68, 0, 0, 0, 0, 0, 0, 0, 0),
                (-47984, -50200, -67512, -4428, 36, -108, 7272, 0, 0, 0, 0, 0, 0, 0, 0),
                (-91972, 100, -708, -28, -164, -20, 84, 0, 0, 0, 0, 0, 0, 0, 0),
                (852, 28, 15760, -1700, 2640, 2644, -460, 0, 0, 0, 0, 0, 0, 0, 0),
                (-668, -11728, -1548, 332, 1724, -3892, 92868, 0, 0, 0, 0, 0, 0, 0, 0),
                (28, -8932, -59664, 12, 4628, -74200, -76, 0, 0, 0, 0, 0, 0, 0, 0),
                (1396, 1260, -76, -1868, 85356, -6372, 12, 0, 0, 0, 0, 0, 0, 0, 0)
                );
    constant children_left : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 13, 9, 11, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1),
                (1, 3, 5, 7, 9, 11, 13, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant children_right : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 14, 10, 12, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1),
                (2, 4, 6, 8, 10, 12, 14, -1, -1, -1, -1, -1, -1, -1, -1)
                );
    constant value_int : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 0, 0, 0, 0, 0, 0, -4, 4, -1, -5, 0, -4, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, 1, -4, -3, -4, -4, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 2, 0, -4, -1, -3, 1, -3),
                (0, 0, 0, 0, 0, 0, 0, -3, 0, -2, -4, 2, -2, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, -3, 0, -2, 0, 1, -2, -3, -1),
                (0, 0, 0, 0, 0, 0, 0, 2, -2, -2, 1, -3, -2, 0, 2),
                (0, 0, 0, 0, 0, 0, 0, -2, -4, 2, -3, 0, -2, -3, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, -1, -3, 1, -1, -1, 3),
                (0, 0, 0, 0, 0, 0, 0, -2, -1, 1, -1, -3, 1, 3, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, -3, 1, 0, -3, -2, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -1, 1, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -2, 1, -1, -2, -1, -3, 1),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, -3, -1, -2, 1, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, -3, 2, -2, 0, -2, 1, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -2, -1, -2, 0, 2, -2),
                (0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 1, -3, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, 1, 0, -2, -1, 0, 3),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, -3, 1, 2, -1, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, 1, -1, -2, 0, 1, 3),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, 1, -2, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -3, -1, 1, -1, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, -3, -1, 0, -2, 1, 1, -2, 3),
                (0, 0, 0, 0, 0, 0, 0, -4, -2, -2, 0, -1, 0, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 1, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, 0, -2, 1, -1, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, -1, 1, -1, 0, 1, -3, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -2, 1, -1, 0, -3, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, -2, -1, -2, 0, 0, 0, -2, -1),
                (0, 0, 0, 0, 0, 0, 0, 1, -2, -1, 0, -1, 2, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, -1, -3, 0, -2, -1, 1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 4, 1, -1, 0, -1, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 1, 0, -1, 2),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, -3, -1, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, 0, -1, -2, -1, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 0, -2, 0, -2, -1),
                (0, 0, 0, 0, 0, 0, 0, 13, 3, -1, 0, 1, -1, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, -2, -2, 4),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -3, -1, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, -4, -1, 0, 0, -2, 0, 1, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, -2, -4, -3, -1, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, -2, 0, -1, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1, -5, 2, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -2, -2, 1),
                (0, 0, 0, 0, 0, 0, 0, 2, -21, -1, 2, -2, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, -2, 0, -1, -3, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -3, -1, -2, 0, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -3, 0, -1, 0, -1, 1, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -3, 0, -2, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -2, -1, 1, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 1, 1, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, -1, 1, -1, 0, -1, 1),
                (0, 0, 0, 0, 0, 0, 0, 5, -2, 0, 0, -3, 1, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, 3, -1, -2, -3, -2, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, 1, -2, 0, -3, 1, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, -2, 1, 0, 0, -1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, -3, 0, 0, 1, 0, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, -2, 1, -3, -2, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, 1, -1, -2, 0, -2, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -4, -3, 2, 0, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, 0, 0, -2, 1, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, -1, 0, 0, -1, 2, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, -2, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, -14, 1, -1, 0, -3, 0, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, -1, -2, 1, -2),
                (0, 0, 0, 0, 0, 0, 0, 0, -3, 9, 2, 0, 0, -2, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, -4, 0, 0, -2, 1, 1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -3, -2, -4, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 3, 14, -1, 0, 0, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 0, -3, -1, -1, -3, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 6, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -2, -1, -3, -1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -3, -1, -3, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -3, 0, -1, -4, -1, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, 1, 0, 1, 0, 0, -1, 0),
                (0, 0, 0, 0, 32, 0, 0, 1, 3, 0, -2, 0, 0, 32, 32),
                (0, 0, 0, 0, 0, 0, 0, 0, -2, 0, 1, 0, -1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 8, -3, 0, 0, 0, -1, -3),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, -1, 0, 1, 0),
                (0, 0, 0, 0, 0, 0, 0, 2, -1, -2, -1, 0, -2, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 5, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 1, -1, -1, 0, 0, -2),
                (0, 0, 0, 0, 0, 0, 0, -2, 2, 0, -2, 0, 0, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, -2, 2, -1, 4, -1),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -2, 7, -1, -2, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -2, -1, 3, -1, 0, 0, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 0, -3, 0, 0, -2, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, 1, -1, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, 6, 2, -2, 0, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, -1, -3, 0, -3, -6, 0, 2),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -4, 0, -1, 1, -2, -1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 0, 0, -1, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, -1, 2, 0, -1, 0, 0, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 1, -2, 0, 1, 0, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -3, 0, 1, -1, 0, -1),
                (0, 0, 0, 0, 0, 0, 0, -1, 1, -3, -1, 1, -3, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 1, 0, -1, 0, 0, 0, 2, 0),
                (0, 0, 0, 0, 0, 0, 0, 7, -2, 0, 0, -2, 6, 7, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 3, -2, 1, 0, -1, 0, 1),
                (0, 0, 0, 0, 0, 0, 0, 2, 10, -1, 0, 0, -2, 0, 0),
                (0, 0, 0, 0, 0, 0, 0, 0, 0, -1, 1, 3, 0, -2, 0)
                );
    constant parent : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 5, 5, 6, 6, 4, 4),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6),
                (-1, 0, 0, 1, 1, 2, 2, 3, 3, 4, 4, 5, 5, 6, 6)
                );
    constant depth : intArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := ((0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3),
                (0, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3)
                );
    constant iLeaf : intArray2D(nTrees-1 downto 0)(nLeaves-1 downto 0) := ((7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14),
                (7, 8, 9, 10, 11, 12, 13, 14)
                );
    constant value : tyArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_tyArray2D(value_int);
      constant threshold : txArray2D(nTrees-1 downto 0)(nNodes-1 downto 0) := to_txArray2D(threshold_int);
end Arrays0;